/sos/cache/7/Projects-BIN.cac/CCE7502/FILES/logic#lib#lef#pll#lef_128_82