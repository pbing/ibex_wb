/sos/cache/7/Projects-BIN.cac/CCE7502/FILES/logic#lib#lef#xtal#lef_129_83